let x = fun y -> y + 1 in
(x 1)